module processor();
/**inputs : instrucction memory, clock, readDate, */
/*outputs: dataAddress, readData2, */

endmodule